magic
tech sky130A
magscale 1 2
timestamp 1669849200
<< checkpaint >>
rect 0 0 2520 3520
<< locali >>
rect 432 850 600 910
rect 600 586 864 646
rect 600 586 660 910
rect 324 146 540 206
rect 324 498 540 558
rect 756 938 972 998
rect 2412 132 2628 220
rect -108 132 108 220
<< m3 >>
rect 1548 0 1748 3520
rect 756 0 956 3520
rect 1548 0 1748 3520
rect 756 0 956 3520
use SUNTRB_NDX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2520 704
use SUNTRB_IVX8_CV XA2
transform 1 0 0 0 1 704
box 0 704 2520 3520
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 756 938 972 998 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 4 nsew
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 5 nsew
flabel m3 s 1548 0 1748 3520 0 FreeSans 400 0 0 0 AVDD
port 6 nsew
flabel m3 s 756 0 956 3520 0 FreeSans 400 0 0 0 AVSS
port 7 nsew
<< end >>
