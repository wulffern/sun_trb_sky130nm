magic
tech sky130B
magscale 1 2
timestamp 1709161200
<< checkpaint >>
rect 0 0 2520 704
<< locali >>
rect 834 234 894 470
rect 1626 234 1686 470
rect 864 586 1032 646
rect 1032 586 1656 646
rect 1032 586 1092 646
rect 324 146 540 206
rect 1980 498 2196 558
rect 324 498 540 558
rect 756 586 972 646
rect 2412 132 2628 220
rect -108 132 108 220
<< poly >>
rect 324 158 2196 194
<< m3 >>
rect 1548 0 1748 704
rect 756 0 956 704
rect 1548 0 1748 704
rect 756 0 956 704
use SUNTRB_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTRB_NCHDL MN1 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTRB_PCHDL MP0 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTRB_PCHDL MP1 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTRB_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use SUNTRB_cut_M1M4_2x1 xcut1 
transform 1 0 756 0 1 58
box 756 58 956 134
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 1980 498 2196 558 0 FreeSans 400 0 0 0 CN
port 3 nsew signal bidirectional
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 C
port 2 nsew signal bidirectional
flabel locali s 756 586 972 646 0 FreeSans 400 0 0 0 Y
port 4 nsew signal bidirectional
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 5 nsew signal bidirectional
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 6 nsew signal bidirectional
flabel m3 s 1548 0 1748 704 0 FreeSans 400 0 0 0 AVDD
port 7 nsew signal bidirectional
flabel m3 s 756 0 956 704 0 FreeSans 400 0 0 0 AVSS
port 8 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 704
<< end >>
